`timescale 1ns/1ps
module egakzxppxv(in0, in2, clock_1, out51);
  wire _0090_;
  reg _0200_ = 1;
  reg [10:0] _0216_ = 1;
  wire [11:0] _0258_;
  reg [22:0] _0274_ = 1;
  wire [16:0] _0539_;
  input clock_1;
  input [23:11] in0;
  input [27:8] in2;
  wire [21:5] out21;
  output out51;
  reg [24:15] reg_18 = 10'h000;
  assign _0104_ = ! _0509_;
  assign _0201_ = _0258_ > 12'hab7;
  assign _0204_ = 7'h7f <= _0104_;
  assign _0258_ = 3'h3 ||  _0274_;
  always @(negedge clock_1, posedge in0)
    if (_0090_) reg_18 <= 10'h09d;
  assign _0412_ = | reg_18[19:18];
  assign _0413_ = | _0537_;
  assign _0537_ = in2[11] ?  11'h03e : _0216_;
  assign _0538_ = _0412_ ?  out21 : _0201_;
  assign _0539_ = _0413_ ?  _0538_ : 17'h00570;
  assign out21 = _0204_;
  assign out51 = _0539_[0];
  assign _0509_ = _0200_;
endmodule
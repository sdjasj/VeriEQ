`timescale 1ns/1ps
module itmozsmldb (in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, clock_0, clock_1, clock_2, clock_3, clock_4, clock_5, clock_6, clock_7, clock_8, clock_9, clock_10, clock_11, clock_12, clock_13, clock_14, clock_15, clock_16, clock_17, clock_18, clock_19, out0, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12, out13, out14, out15, out16, out17, out18, out19 );

input wire in0;
input wire [28:18] in1;
input wire [31:15] in2;
input wire [1:0] in3;
input wire in4;
input wire [30:24] in5;
input wire [19:9] in6;
input wire [11:8] in7;
input wire [10:2] in8;
input wire [10:8] in9;
input wire [19:7] in10;
input wire [21:15] in11;
input wire [18:14] in12;
input wire [12:5] in13;
input wire [24:13] in14;
input wire in15;
input wire [12:4] in16;
input wire [20:10] in17;
input wire [35:15] in18;
input wire [10:5] in19;
wire wire_0;
wire wire_1;
wire wire_2;
wire [15:11] wire_3;
wire [7:2] wire_4;
wire [2:1] wire_5;
wire [31:6] wire_6;
wire [2:2] wire_7;
wire [21:16] wire_8;
wire wire_9;
reg [27:6] reg_0;
reg reg_1;
reg [1:0] reg_2;
reg [17:2] reg_3;
reg reg_4;
reg reg_5;
reg [23:19] reg_6;
reg reg_7;
reg reg_8;
reg [17:2] reg_9;
reg reg_10;
reg [30:10] reg_11;
reg reg_12;
reg [8:2] reg_13;
reg [3:3] reg_14;
reg [16:8] reg_15;
reg reg_16;
reg reg_17;
reg [25:16] reg_18;
reg [26:18] reg_19;
reg [26:1] reg_20;
reg reg_21;
reg reg_22;
reg [8:6] reg_23;
reg [31:19] reg_24;
reg [3:1] reg_25;
reg [1:1] reg_26;
reg [30:15] reg_27;
reg reg_28;
reg [33:13] reg_29;
reg [7:7] reg_30;
reg [6:3] reg_31;
reg reg_32;
reg [24:5] reg_33;
reg reg_34;
reg reg_35;
reg [16:6] reg_36;
reg reg_37;
reg [18:14] reg_38;
reg [23:3] reg_39;
reg [25:7] reg_40;
reg [0:0] reg_41;
reg reg_42;
reg [27:15] reg_43;
reg [23:11] reg_44;
reg [26:20] reg_45;
reg [27:13] reg_46;
reg reg_47;
reg reg_48;
reg [14:9] reg_49;
reg [25:22] reg_50;
output wire out0;
output wire out1;
output wire [11:3] out2;
output wire [8:1] out3;
output wire [23:9] out4;
output wire [32:20] out5;
output wire [0:0] out6;
output wire [4:4] out7;
output wire [34:8] out8;
output wire [35:16] out9;
output wire [30:18] out10;
output wire out11;
output wire out12;
output wire [17:0] out13;
output wire [19:8] out14;
output wire [7:6] out15;
output wire [17:13] out16;
output wire [10:0] out17;
output wire out18;
output wire out19;
input clock_0;
wire clock_0;
input clock_1;
wire clock_1;
input clock_2;
wire clock_2;
input clock_3;
wire clock_3;
input clock_4;
wire clock_4;
input clock_5;
wire clock_5;
input clock_6;
wire clock_6;
input clock_7;
wire clock_7;
input clock_8;
wire clock_8;
input clock_9;
wire clock_9;
input clock_10;
wire clock_10;
input clock_11;
wire clock_11;
input clock_12;
wire clock_12;
input clock_13;
wire clock_13;
input clock_14;
wire clock_14;
input clock_15;
wire clock_15;
input clock_16;
wire clock_16;
input clock_17;
wire clock_17;
input clock_18;
wire clock_18;
input clock_19;
wire clock_19;


	initial begin
		#1;
		    reg_0 = 0;
    reg_1 = 0;
    reg_2 = 0;
    reg_3 = 0;
    reg_4 = 0;
    reg_5 = 0;
    reg_6 = 0;
    reg_7 = 0;
    reg_8 = 0;
    reg_9 = 0;
    reg_10 = 0;
    reg_11 = 0;
    reg_12 = 0;
    reg_13 = 0;
    reg_14 = 0;
    reg_15 = 0;
    reg_16 = 0;
    reg_17 = 0;
    reg_18 = 0;
    reg_19 = 0;
    reg_20 = 0;
    reg_21 = 0;
    reg_22 = 0;
    reg_23 = 0;
    reg_24 = 0;
    reg_25 = 0;
    reg_26 = 0;
    reg_27 = 0;
    reg_28 = 0;
    reg_29 = 0;
    reg_30 = 0;
    reg_31 = 0;
    reg_32 = 0;
    reg_33 = 0;
    reg_34 = 0;
    reg_35 = 0;
    reg_36 = 0;
    reg_37 = 0;
    reg_38 = 0;
    reg_39 = 0;
    reg_40 = 0;
    reg_41 = 0;
    reg_42 = 0;
    reg_43 = 0;
    reg_44 = 0;
    reg_45 = 0;
    reg_46 = 0;
    reg_47 = 0;
    reg_48 = 0;
    reg_49 = 0;
    reg_50 = 0;

	end
    assign wire_0 = (in4 ^ in4) ? (12'o7634 || !(in2[24:24]) ? 3'b10 : (9'd386 || 8'hb3)) ? 7'o127 ? in1 : 9'd497 ? (in11[17:17] & 4'h09) : 2'o03 ? 2'h2 : in3 ? in4 ? (5'b01 >> in16[9:8]) : -(in19[6:6]) : in11[15:15] : ~(9'd257) : -((in9[8:8] && 4'ha)) ? (in17[18:18] << in12[16:16]) : in11[19:19] ? in14[17:17] : in8[5:4];
    assign wire_1 = in11[17:17];
    assign wire_2 = 4'ha;
    assign wire_3 = 6'b110;
    assign wire_4 = in0;
    assign wire_5 = in1[26:26] ? wire_1 : 10'd783;
    assign wire_6 = 7'h5a ? (!(12'hc0a) && ((12'hb40 * 12'o7223) % ({1'b1, -(in18[16:16])})) ? ~(wire_2) ? 6'o44 : 13'b100000001 ? in16[4:4] : in8[3:3] : 9'o775) : in9;
    assign wire_7 = in18[29:18];
    assign wire_8 = -(~(wire_6[17:16]));
    assign wire_9 = 6'o62;
    assign out0 = 12'o7167;
    assign out1 = reg_20;
    assign out2 = 6'h27;
    assign out3 = 8'b00001 ? ((in4 ^ 10'd881) || (3'o6 >= 3'h6)) : 5'b0 ? 1'o1 ? 10'o1733 : (-(reg_46[13:13]) ? reg_41[0:0] : 9'b100110 - 8'b11100 ? in10[7:7] ? reg_14 : reg_16 : !(reg_28)) : ((wire_3[12:12] * 12'hd9d) ? !(9'b1000000) : 3'h7 < (8'o363 || 9'o441 ? in18[27:27] : out0)) ? in1[28:28] : reg_33[15:14];
    assign out4 = -((-(!(reg_9[6:6])) ? 8'd217 : 10'd830 ? 7'b11110 : in9[9:9] ? reg_33[12:10] : reg_16 + ((reg_0[20:20] && 6'b000101) ? 5'o024 : ~(in2[22:20]) ~^ 4'ha ? 6'b1 ? reg_43[24:23] : wire_7[2:2] : ~(wire_2))));
    assign out5 = wire_6[9:7];
    assign out6 = 10'd874;
    assign out7 = ~(3'o007 ? (out2 ? 5'd22 ? 8'hf6 : wire_4[2:2] : wire_0 << reg_3[11:11]) : ~(7'd118) ? 9'd273 : (10'd629 ^ in4 ? 10'd801 : 4'hd));
    assign out8 = (((12'o4014 < reg_31[6:6]) || reg_43[16:16]) % ({1'b1, -((10'd685 && 3'o5))})) ? (!(out6) > 2'o2) : 11'b100001000 ? !(reg_12 ? ~(reg_33[11:11]) : (wire_8[16:16] <= 11'o3154) ? !((10'd606 == wire_7[2:2])) : 10'd687 ? reg_35 : 10'b1010110 ? (13'b01011001 <= in13[12:11]) : 8'he9) : reg_47;
    assign out9 = -(wire_6[20:20]);
    assign out10 = !(((reg_30[7:7] && reg_36) ? ~(reg_24[20:20]) : -(8'd199) ? ~(reg_24[28:28]) : (11'o3056 >= (6'b11011 == wire_4[5:5])) * (5'o33 | !(reg_6) ? (8'd228 != reg_18[18:18]) : 2'b0)));
    assign out11 = 9'd447 ? -(reg_14) : reg_14[3:3];
    assign out12 = (reg_35 << ((-(in15) % ({1'b1, !(wire_5[1:1])})) / ({1'b1, 4'hd})) ? !((reg_0[21:13] && 7'h56)) ? 4'b11 : ~(reg_6[21:21] ? 9'd264 : reg_48) : 10'd749);
    assign out13 = (reg_42 & ~(in10[15:15])) ? 7'd87 : !((!(wire_6[8:8]) | 10'd740)) ? reg_13[7:7] ? ~(8'd156) : ((reg_27[26:25] & 10'd918) & reg_36[9:8]) : reg_41;
    assign out14 = 6'o056;
    assign out15 = 3'o5;
    assign out16 = ((-(7'o116) + in7) > 2'o3 ? !(reg_35) : (out2[7:6] && reg_40[11:8]) ? -(10'd583 ? reg_11[21:18] : 9'h181) : !(in13[5:5]) ? (out6[0:0] << 7'd101) : out10[21:20] ? reg_40[9:9] : reg_28 ? out3[1:1] : !(~(reg_18)) ? (out15[7:7] ? reg_27[15:15] : reg_2 && reg_15[11:9]) : (!(in16) * 9'd503 ? 10'd758 : 3'b00));
    assign out17 = 12'he1c;
    assign out18 = !(!(4'he));
    assign out19 = (-((in17[16:16] >> reg_3[2:2]) ? 9'd256 : reg_23[6:6]) >= !(wire_5[2:2] ? (9'd490 ? reg_0[12:10] : in15 < -(wire_1)) : 1'o0));
always @(negedge clock_15 or posedge clock_2 or negedge clock_18 or negedge clock_9 or negedge clock_8 or posedge clock_10 or negedge clock_3 or negedge clock_17 or posedge clock_11 or negedge clock_5 or posedge clock_16 or negedge clock_1 or posedge clock_6 or posedge clock_12) begin
  if (clock_12) begin
    reg_0 <= 569;
    reg_1 <= 569;
    reg_2 <= 569;
    reg_3 <= 569;
    reg_4 <= 569;
    reg_5 <= 569;
    reg_6 <= 569;
    reg_7 <= 569;
    reg_8 <= 569;
    reg_9 <= 569;
    reg_10 <= 569;
    reg_11 <= 569;
    reg_12 <= 569;
    reg_13 <= 569;
    reg_14 <= 569;
    reg_15 <= 569;
    reg_16 <= 569;
    reg_17 <= 569;
    reg_18 <= 569;
    reg_19 <= 569;
    reg_20 <= 569;
    reg_21 <= 569;
    reg_22 <= 569;
    reg_23 <= 569;
    reg_24 <= 569;
    reg_25 <= 569;
  end else begin
  if (in8[2:2]) begin
  reg_0[24:18] <= wire_8[16:16];
  reg_1 <= (in6 ? 8'hd2 : !(wire_7[2:2] ? in12[15:15] : in8[4:4]) ? in0 : 7'b1100101 == 8'b11111);
end else begin
  reg_2[1:0] <= wire_7[2:2];
  reg_3[6:5] <= !(~(in4) ? (8'h8f ? 11'h5c3 : in0 ? wire_2 : wire_8[18:18] >= -(in15)) : (in2[21:21] - (wire_1 >> in14[20:19])));
end
  case (7'b000111)
  10'd633: begin
    reg_4 <= (13'b0111001010 % ({1'b1, 10'd626}));
    reg_5 <= ((-(~((9'd355 >> in10))) != -(in9[10:10]) ? !(wire_7[2:2]) : wire_1 ? (5'b010 && 10'd600) ? (wire_0 >> in1[19:19]) : in19[5:5] ? in6 : in10[7:7] : ~((10'd862 | 5'b110))) && (wire_7 ~^ 10'd830));
    reg_6[19:19] <= ~(((wire_8[16:16] << in18[16:16]) % ({1'b1, 4'o16})) ? 3'o5 : ((~(in6[12:12]) * !(10'd747)) ^ wire_0));
  end
  11'b100100100: begin
    reg_7 <= ((in13[5:5] >> (wire_3[13:13] / ({1'b1, ~(in2[18:17])}))) <= 4'hd);
    reg_8 <= 2'o3 ? 1'o0 : in1[27:27];
  end
  default: begin
    reg_9[10:4] <= 10'd599 ? ~((!((in5[25:25] && wire_6[11:11])) > in13)) : wire_7[2:2];
  end
endcase
  if (wire_0) begin
  reg_10 <= 1'o1;
  reg_11[20:20] <= -(-(in13[8:7]) ? 4'he : -(wire_0) ? -(in9[9:8]) : !((5'd18 * 8'd239)) ? in8[10:10] ? -(in2[26:25]) : !(in5[24:24]) ? (in5[24:24] << 8'h96) : 4'd12 : 5'b0100);
  reg_12 <= in14[19:19] ? ((~(4'hc) * in9[9:8]) & 6'b0000) : in9;
end else begin
  reg_13[4:3] <= (in5[26:26] - (wire_6[17:17] ? (4'o13 ^ in9[9:9]) ? 6'b0000 ? 9'd376 : 10'd544 : ~(8'd189) : in17[16:16] ~^ -(wire_5[1:1] ? in17[17:15] : !(10'd989))));
  reg_14[3:3] <= (!(wire_1) != 12'hac0);
  reg_15[11:9] <= in15;
end
  case (14'b1001110111)
  8'd178: begin
    reg_16 <= (-((in8[7:7] ? 10'b101110 : wire_6[23:21] < 9'o661)) < 8'b11100 ? ~(9'd345) : 9'o747) ? -(4'b01 ? 4'hb : 10'b0111111010 ? (9'b0110 >> 10'd938) ? 12'o5126 : in1[20:19] : ~((9'd350 / ({1'b1, in7[10:9]})))) : 7'h7c;
  end
  5'o36: begin
    reg_17 <= ~((wire_9 << 2'b0 ? (9'd341 + in1[23:23]) : 9'b1111000) ? (~(8'hbe) | in17[12:12]) ? (in2[16:16] ? wire_5[1:1] : in5[27:27] - !(8'hf6)) : in8[5:5] ? in6[11:11] : 11'b0000111 : in3[0:0]);
    reg_18[19:18] <= (~((wire_9 - 12'b0010111)) / ({1'b1, in1})) ? in11 ? (9'o614 > wire_5[1:1]) : (in15 + (in12[14:14] ~^ 6'o61)) : in8[4:4] ? (in9 * (-(5'o37) ? (in17[20:20] << in18[17:17]) : 6'o062 << (in10 ~^ in11))) : 8'o0216;
  end
  12'o5132: begin
    reg_19[26:18] <= 2'o3;
    reg_20[18:7] <= in19[6:6];
  end
  8'd203: begin
    reg_21 <= 3'b101 ? 6'o71 : (((8'b1010000 && 6'd61) | (in17 / ({1'b1, 12'b00100111}))) == 10'd870 ? 10'b0110101 ? 8'h83 : wire_0 : !(8'h8c)) ? 8'd234 : -(-(9'o712) ? 9'd326 ? 12'b1100010 : in12[14:14] : in0);
  end
  default: begin
    reg_22 <= in16;
    reg_23[8:6] <= 10'd980;
    reg_24[29:21] <= in6[9:9];
  end
endcase
  reg_25[2:2] <= ~(12'o5231);
  end
end
always @(posedge clock_3 or posedge clock_12 or negedge clock_4 or posedge clock_11 or posedge clock_14 or negedge clock_1 or negedge clock_6 or negedge clock_19 or negedge clock_18 or negedge clock_16 or negedge clock_15 or posedge clock_2 or negedge clock_17 or posedge clock_0 or posedge clock_10 or negedge clock_13 or negedge clock_9 or posedge clock_5) begin
  if (clock_5) begin
    reg_26 <= 721;
    reg_27 <= 721;
    reg_28 <= 721;
    reg_29 <= 721;
    reg_30 <= 721;
    reg_31 <= 721;
    reg_32 <= 721;
    reg_33 <= 721;
    reg_34 <= 721;
  end else begin
  reg_26[1:1] <= (10'b0000100101 >= (2'o3 < wire_0)) ? wire_6[23:20] : (6'd50 ? 1'h0 : 12'o6067 > !(12'hcfe)) ? 9'd335 ? reg_23 : in7 ? (12'o7735 && in1[25:25]) : in12[15:14] : -(in13) ? reg_11[17:15] ? wire_5[1:1] ? 10'd788 : wire_2 : 7'd111 ? reg_8 : (12'o6070 ? in7[9:8] : 10'd782 >> reg_6[20:20] ? 8'b00001100 : 8'hb1) : wire_8[16:16] ? 10'd603 : 10'd636 ? 12'hba4 : 10'd691 ? in6[10:10] : in5[24:24];
  if ((~(((!(wire_5[1:1]) ~^ 4'hf ? in14[21:20] : in3[0:0]) ~^ 10'b001011101)) >= 4'b010)) begin
  reg_27[22:18] <= 8'b1101011;
  reg_28 <= 6'b1;
  reg_29[22:15] <= in3[0:0];
end else begin
  reg_30[7:7] <= 7'd112;
  reg_31[5:4] <= -(4'b100);
end
  reg_32 <= reg_2[1:0] ? (!(in17[19:17]) | reg_13[6:6] ? reg_19 : reg_17) : ~(!(!(-(1'h1))));
  reg_33[18:13] <= wire_2;
  reg_34 <= !((in12[14:14] >= ((wire_1 + 6'o76) / ({1'b1, (1'b0 > 12'o5423)})))) ? 5'b10 : 8'h90;
  end
end
always @(posedge clock_17 or negedge clock_15 or negedge clock_0 or posedge clock_12 or posedge clock_19 or posedge clock_11 or negedge clock_6 or negedge clock_10 or negedge clock_14 or negedge clock_5 or posedge clock_7 or negedge clock_13 or posedge clock_1 or posedge clock_3 or negedge clock_16 or negedge clock_4 or posedge clock_18) begin
  if (clock_18) begin
    reg_35 <= 545;
    reg_36 <= 545;
    reg_37 <= 545;
    reg_38 <= 545;
    reg_39 <= 545;
    reg_40 <= 545;
    reg_41 <= 545;
    reg_42 <= 545;
    reg_43 <= 545;
    reg_44 <= 545;
    reg_45 <= 545;
    reg_46 <= 545;
    reg_47 <= 545;
    reg_48 <= 545;
    reg_49 <= 545;
    reg_50 <= 545;
  end else begin
  reg_35 <= (reg_3[3:2] == reg_7);
  reg_36[10:6] <= in1[26:22];
  case (7'b000)
  13'b11100110: begin
    reg_37 <= 9'b001111;
    reg_38[18:18] <= in0;
  end
  4'hb: begin
    reg_39[3:3] <= (-(in6[9:9]) < ((reg_3[7:6] >> in6[9:9] ? reg_18[18:18] : reg_0[22:19]) ? 10'd514 : wire_1 << reg_12));
    reg_40[22:18] <= reg_7;
  end
  8'd137: begin
    reg_41[0:0] <= ~(reg_26);
    reg_42 <= -(reg_7);
  end
  default: begin
    reg_43[25:23] <= wire_8[18:18];
    reg_44[19:17] <= !(9'o410);
    reg_45[24:20] <= 5'o23;
  end
endcase
  case (reg_14[3:3])
  10'd516: begin
    reg_46[24:22] <= 3'o6;
  end
  8'he7: begin
    reg_47 <= -(-(3'o6 ? 11'h64f : ((in0 & 3'o05) % ({1'b1, 8'd166 ? wire_8[18:17] : 11'b1100011010}))));
  end
  default: begin
    reg_48 <= ~(!(3'o5));
    reg_49[12:10] <= (in18[26:26] >= ~(~(13'b1101010111)) ? (3'h4 == ~(3'h7)) : reg_19[23:23] ? (reg_30[7:7] / ({1'b1, (6'h38 ? 7'd95 : 10'd791 <= in2[15:15])})) : (reg_18 || 7'b110101) ? in5[28:28] ? reg_16 : wire_3 : 4'h8 ? reg_25[1:1] : 6'o45 ? reg_31 : ~(-(6'b1011)));
  end
endcase
  reg_50[24:24] <= in13[6:6];
  end
end
endmodule

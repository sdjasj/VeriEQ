module top(input a, output b);
  begin
    
  end
endmodule